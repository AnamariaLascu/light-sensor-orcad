** Profile: "SCHEMATIC1-sim_tranzitoriu"  [ c:\cadence\lascuanamaria_orcad\proiect_cad-PSpiceFiles\SCHEMATIC1\sim_tranzitoriu.sim ] 

** Creating circuit file "sim_tranzitoriu.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../proiect_cad-pspicefiles/verde.lib" 
.LIB "../../../proiect_cad-pspicefiles/rosu.lib" 
.LIB "../../../proiect_cad-pspicefiles/portocaliu.lib" 
.LIB "../../../proiect_cad-pspicefiles/galben.lib" 
.LIB "../../../proiect_cad-pspicefiles/albastru.lib" 
* From [PSPICE NETLIST] section of C:\Users\Ana\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "C:\Cadence\LascuAnamaria_orCAD\proiect1-PSpiceFiles\blue.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 200us 0 2u 
.STEP LIN PARAM senzor 25k 40k 1k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
